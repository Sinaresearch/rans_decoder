
// tables from the C code that go with the algorithm.  These tables must be 
// regenerated for every input file!  They are unique to each encoding.
// Do not change the input file without making new tables!


`timescale 1ns / 1ns
module ANSTables(
input [7:0]divider_index,
input [8:0]slot_adjust_index,
input [8:0]sym_id_index,
input [8:0]slot_freqs_index,
output wire [31:0]dividerQ,
output wire [31:0]slot_adjustQ,
output wire [31:0]sym_idQ,
output wire [31:0]slot_freqsQ
);

parameter NSYM = 256;
parameter WORD_WIDTH = 32;
wire [WORD_WIDTH * NSYM-1:0]divider;
wire [WORD_WIDTH * NSYM * 2-1:0]slot_adjust;
wire [WORD_WIDTH * NSYM * 2-1:0]sym_id;
wire [WORD_WIDTH * NSYM * 2-1:0]slot_freqs;


// perform table lookup given index into table.
assign dividerQ = divider[((NSYM - divider_index-1)*WORD_WIDTH)+:WORD_WIDTH];
assign slot_adjustQ = slot_adjust[((NSYM*2-slot_adjust_index-1)*WORD_WIDTH)+:WORD_WIDTH];
assign sym_idQ = sym_id[((NSYM*2-sym_id_index-1)*WORD_WIDTH)+:WORD_WIDTH];
assign slot_freqsQ = slot_freqs[((NSYM*2-slot_freqs_index-1)*WORD_WIDTH)+:WORD_WIDTH];



// Start of Computer Generated tables:

assign divider = {
32'h00000000, 32'h00000100, 32'h00000200, 32'h00000300, 32'h00000400, 32'h00000500, 32'h00000600, 32'h00000700, 32'h00000800, 32'h00000900, 32'h00000a39, 32'h00000b00, 32'h00000c00, 32'h00000d00, 32'h00000e00, 32'h00000f00, 
32'h00001000, 32'h00001100, 32'h00001200, 32'h00001300, 32'h00001400, 32'h00001500, 32'h00001600, 32'h00001700, 32'h00001800, 32'h00001900, 32'h00001a00, 32'h00001b00, 32'h00001c00, 32'h00001d00, 32'h00001e00, 32'h00001f00, 
32'h00002093, 32'h00002100, 32'h00002200, 32'h00002300, 32'h00002400, 32'h00002500, 32'h00002600, 32'h00002700, 32'h00002800, 32'h00002900, 32'h00002a00, 32'h00002b00, 32'h00002c76, 32'h00002d05, 32'h00002ec7, 32'h00002f00, 
32'h00003000, 32'h00003100, 32'h00003200, 32'h00003300, 32'h00003400, 32'h00003500, 32'h00003600, 32'h00003700, 32'h00003800, 32'h00003900, 32'h00003a00, 32'h00003b00, 32'h00003c00, 32'h00003d00, 32'h00003e00, 32'h00003f00, 
32'h00004000, 32'h0000415b, 32'h00004200, 32'h0000438e, 32'h00004456, 32'h000045e4, 32'h00004655, 32'h00004700, 32'h000048c7, 32'h0000491d, 32'h00004a00, 32'h00004bc7, 32'h00004c00, 32'h00004dc7, 32'h00004ee4, 32'h00004f5c, 
32'h000050c7, 32'h00005100, 32'h0000528f, 32'h000053c7, 32'h0000543a, 32'h00005500, 32'h00005600, 32'h000057c7, 32'h00005800, 32'h00005900, 32'h00005a00, 32'h00005b00, 32'h00005c00, 32'h00005d00, 32'h00005e00, 32'h00005f00, 
32'h00006000, 32'h000061d1, 32'h00006200, 32'h00006372, 32'h00006460, 32'h0000657f, 32'h000066d5, 32'h000067f2, 32'h000068d7, 32'h00006967, 32'h00006a00, 32'h00006b4b, 32'h00006c2f, 32'h00006dda, 32'h00006ef8, 32'h00006fc0, 
32'h000070a4, 32'h00007100, 32'h000072a6, 32'h00007319, 32'h0000748c, 32'h000075c6, 32'h000076c7, 32'h000077e3, 32'h000078c7, 32'h00007a00, 32'h00007a00, 32'h00007b00, 32'h00007c00, 32'h00007d00, 32'h00007e00, 32'h00007f00, 
32'h00008000, 32'h00008100, 32'h00008200, 32'h00008300, 32'h00008400, 32'h00008500, 32'h00008600, 32'h00008700, 32'h00008800, 32'h00008900, 32'h00008a00, 32'h00008b00, 32'h00008c00, 32'h00008d00, 32'h00008e00, 32'h00008f00, 
32'h00009000, 32'h00009100, 32'h00009200, 32'h00009300, 32'h00009400, 32'h00009500, 32'h00009600, 32'h00009700, 32'h00009800, 32'h00009900, 32'h00009a00, 32'h00009b00, 32'h00009c00, 32'h00009d00, 32'h00009e00, 32'h00009f00, 
32'h0000a000, 32'h0000a100, 32'h0000a200, 32'h0000a300, 32'h0000a400, 32'h0000a500, 32'h0000a600, 32'h0000a700, 32'h0000a800, 32'h0000a900, 32'h0000aa00, 32'h0000ab00, 32'h0000ac00, 32'h0000ad00, 32'h0000ae00, 32'h0000af00, 
32'h0000b000, 32'h0000b100, 32'h0000b200, 32'h0000b300, 32'h0000b400, 32'h0000b500, 32'h0000b600, 32'h0000b700, 32'h0000b800, 32'h0000b900, 32'h0000ba00, 32'h0000bb00, 32'h0000bc00, 32'h0000bd00, 32'h0000be00, 32'h0000bf00, 
32'h0000c000, 32'h0000c100, 32'h0000c200, 32'h0000c300, 32'h0000c400, 32'h0000c500, 32'h0000c600, 32'h0000c700, 32'h0000c800, 32'h0000c900, 32'h0000ca00, 32'h0000cb00, 32'h0000cc00, 32'h0000cd00, 32'h0000ce00, 32'h0000cf00, 
32'h0000d000, 32'h0000d100, 32'h0000d200, 32'h0000d300, 32'h0000d400, 32'h0000d500, 32'h0000d600, 32'h0000d700, 32'h0000d800, 32'h0000d900, 32'h0000da00, 32'h0000db00, 32'h0000dc00, 32'h0000dd00, 32'h0000de00, 32'h0000df00, 
32'h0000e000, 32'h0000e100, 32'h0000e200, 32'h0000e300, 32'h0000e400, 32'h0000e500, 32'h0000e600, 32'h0000e700, 32'h0000e800, 32'h0000e900, 32'h0000ea00, 32'h0000eb00, 32'h0000ec00, 32'h0000ed00, 32'h0000ee00, 32'h0000ef00, 
32'h0000f000, 32'h0000f100, 32'h0000f200, 32'h0000f300, 32'h0000f400, 32'h0000f500, 32'h0000f600, 32'h0000f700, 32'h0000f800, 32'h0000f900, 32'h0000fa00, 32'h0000fb00, 32'h0000fc00, 32'h0000fd00, 32'h0000fe00, 32'h0000ff00 
};

assign slot_adjust={
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000100, 32'h00000000, 32'h00000200, 32'h00000000, 32'h00000300, 32'h00000000, 32'h00000400, 32'h00000000, 32'h00000500, 32'h00000600, 32'h00000600, 32'h00000600, 32'h00000700, 
32'h00000600, 32'h00000800, 32'h00000600, 32'h00000900, 32'h00000639, 32'h00000400, 32'h00000639, 32'h00000b00, 32'h00000639, 32'h00000c00, 32'h00000639, 32'h00000d00, 32'h00000639, 32'h00000e00, 32'h00000639, 32'h00000f00, 
32'h00000639, 32'h00001000, 32'h00000639, 32'h00001100, 32'h00000639, 32'h00001200, 32'h00000639, 32'h00001300, 32'h00000639, 32'h00001400, 32'h00000639, 32'h00001500, 32'h00000639, 32'h00001600, 32'h00000639, 32'h00001700, 
32'h00000639, 32'h00001800, 32'h00000639, 32'h00001900, 32'h00000639, 32'h00001a00, 32'h00000639, 32'h00001b00, 32'h00000639, 32'h00001c00, 32'h00000639, 32'h00001d00, 32'h00000639, 32'h00001e00, 32'h00000639, 32'h00001f00, 
32'h00002093, 32'h00000639, 32'h000006a6, 32'h00002100, 32'h000006a6, 32'h00002200, 32'h000006a6, 32'h00002300, 32'h000006a6, 32'h00002400, 32'h000006a6, 32'h00002500, 32'h000006a6, 32'h00002600, 32'h000006a6, 32'h00002700, 
32'h000006a6, 32'h00002800, 32'h000006a6, 32'h00002900, 32'h000006a6, 32'h00002a00, 32'h000006a6, 32'h00002b00, 32'h00002c76, 32'h00002b93, 32'h00002d05, 32'h00002c76, 32'h00002de4, 32'h00002e00, 32'h00002de4, 32'h00002f00, 
32'h00002de4, 32'h00003000, 32'h00003071, 32'h00003100, 32'h00003105, 32'h00003200, 32'h00003300, 32'h00003300, 32'h00003400, 32'h00003400, 32'h00003400, 32'h00003500, 32'h00003600, 32'h00003600, 32'h00003600, 32'h00003700, 
32'h00003600, 32'h00003800, 32'h00003900, 32'h00003900, 32'h00003900, 32'h00003a00, 32'h00003b00, 32'h00003b00, 32'h00003b00, 32'h00003c00, 32'h00003b00, 32'h00003d00, 32'h00003e00, 32'h00003e00, 32'h00003e00, 32'h00003f00, 
32'h00003e00, 32'h00004000, 32'h0000415b, 32'h00003f05, 32'h0000415b, 32'h00004200, 32'h000041e9, 32'h00004200, 32'h0000423f, 32'h00004200, 32'h000045e4, 32'h00004200, 32'h00004639, 32'h00004400, 32'h00004639, 32'h00004700, 
32'h000048c7, 32'h00004800, 32'h000048e4, 32'h00004600, 32'h000048e4, 32'h00004a00, 32'h00004bc7, 32'h00004b00, 32'h00004bc7, 32'h00004c00, 32'h00004c8e, 32'h00004d00, 32'h00004d72, 32'h00004b00, 32'h00004dce, 32'h00004c3f, 
32'h00004e95, 32'h00005000, 32'h00004e95, 32'h00005100, 32'h00004f24, 32'h00005039, 32'h00004feb, 32'h00005300, 32'h00005025, 32'h000051e4, 32'h00005025, 32'h00005500, 32'h00005025, 32'h00005600, 32'h000050ec, 32'h00005700, 
32'h000050ec, 32'h00005800, 32'h000050ec, 32'h00005900, 32'h000050ec, 32'h00005a00, 32'h00005b00, 32'h00005b00, 32'h00005b00, 32'h00005c00, 32'h00005b00, 32'h00005d00, 32'h00005b00, 32'h00005e00, 32'h00005b00, 32'h00005f00, 
32'h00006000, 32'h00006000, 32'h000060d1, 32'h000056ec, 32'h000060d1, 32'h00006200, 32'h00006143, 32'h00005e00, 32'h00006460, 32'h00006143, 32'h0000657f, 32'h00006460, 32'h000066d5, 32'h0000657f, 32'h000067f2, 32'h000066d5, 
32'h000068d7, 32'h000067f2, 32'h00006967, 32'h000068d7, 32'h000066e3, 32'h00006a00, 32'h00006b4b, 32'h00006a67, 32'h00006c2f, 32'h00006b4b, 32'h00006dda, 32'h00006c2f, 32'h00006ef8, 32'h00006dda, 32'h00006fc0, 32'h00006ef8, 
32'h000070a4, 32'h00006fc0, 32'h00006ce3, 32'h00007100, 32'h000072a6, 32'h000071a4, 32'h00007319, 32'h000072a6, 32'h0000748c, 32'h00007319, 32'h000075c6, 32'h0000748c, 32'h000071aa, 32'h00007600, 32'h000077e3, 32'h000076c6, 
32'h00007371, 32'h00007800, 32'h000079e3, 32'h000078e3, 32'h00007471, 32'h00007a00, 32'h00007471, 32'h00007b00, 32'h00007471, 32'h00007c00, 32'h00007be1, 32'h00007d00, 32'h00007be1, 32'h00007e00, 32'h00007be1, 32'h00007f00, 
32'h00007be1, 32'h00008000, 32'h00007be1, 32'h00008100, 32'h00007be1, 32'h00008200, 32'h00007be1, 32'h00008300, 32'h00007be1, 32'h00008400, 32'h00007be1, 32'h00008500, 32'h00007be1, 32'h00008600, 32'h00007be1, 32'h00008700, 
32'h00007be1, 32'h00008800, 32'h00007be1, 32'h00008900, 32'h00007be1, 32'h00008a00, 32'h00007be1, 32'h00008b00, 32'h00007be1, 32'h00008c00, 32'h00007be1, 32'h00008d00, 32'h00007be1, 32'h00008e00, 32'h00007be1, 32'h00008f00, 
32'h00007be1, 32'h00009000, 32'h00007be1, 32'h00009100, 32'h00007be1, 32'h00009200, 32'h00007be1, 32'h00009300, 32'h000092aa, 32'h00009400, 32'h000093e3, 32'h00009500, 32'h000093e3, 32'h00009600, 32'h0000961b, 32'h00009700, 
32'h0000961b, 32'h00009800, 32'h0000961b, 32'h00009900, 32'h0000961b, 32'h00009a00, 32'h0000961b, 32'h00009b00, 32'h0000961b, 32'h00009c00, 32'h0000961b, 32'h00009d00, 32'h0000961b, 32'h00009e00, 32'h0000961b, 32'h00009f00, 
32'h0000961b, 32'h0000a000, 32'h0000a070, 32'h0000a100, 32'h0000a070, 32'h0000a200, 32'h0000a070, 32'h0000a300, 32'h0000a070, 32'h0000a400, 32'h0000a070, 32'h0000a500, 32'h0000a070, 32'h0000a600, 32'h0000a070, 32'h0000a700, 
32'h0000a070, 32'h0000a800, 32'h0000a070, 32'h0000a900, 32'h0000a070, 32'h0000aa00, 32'h0000a070, 32'h0000ab00, 32'h0000a070, 32'h0000ac00, 32'h0000a070, 32'h0000ad00, 32'h0000a070, 32'h0000ae00, 32'h0000a070, 32'h0000af00, 
32'h0000af1c, 32'h0000b000, 32'h0000af1c, 32'h0000b100, 32'h0000af1c, 32'h0000b200, 32'h0000b21c, 32'h0000b300, 32'h0000b21c, 32'h0000b400, 32'h0000b21c, 32'h0000b500, 32'h0000b455, 32'h0000b600, 32'h0000b455, 32'h0000b700, 
32'h0000b455, 32'h0000b800, 32'h0000b7e2, 32'h0000b900, 32'h0000b7e2, 32'h0000ba00, 32'h0000b7e2, 32'h0000bb00, 32'h0000b7e2, 32'h0000bc00, 32'h0000b7e2, 32'h0000bd00, 32'h0000b7e2, 32'h0000be00, 32'h0000b7e2, 32'h0000bf00, 
32'h0000b7e2, 32'h0000c000, 32'h0000b7e2, 32'h0000c100, 32'h0000b7e2, 32'h0000c200, 32'h0000b7e2, 32'h0000c300, 32'h0000b7e2, 32'h0000c400, 32'h0000b7e2, 32'h0000c500, 32'h0000b7e2, 32'h0000c600, 32'h0000b7e2, 32'h0000c700, 
32'h0000b7e2, 32'h0000c800, 32'h0000c838, 32'h0000c900, 32'h0000c838, 32'h0000ca00, 32'h0000c838, 32'h0000cb00, 32'h0000c838, 32'h0000cc00, 32'h0000c838, 32'h0000cd00, 32'h0000c838, 32'h0000ce00, 32'h0000c838, 32'h0000cf00, 
32'h0000cf1c, 32'h0000d000, 32'h0000cf1c, 32'h0000d100, 32'h0000cf1c, 32'h0000d200, 32'h0000d1fe, 32'h0000d300, 32'h0000d1fe, 32'h0000d400, 32'h0000d1fe, 32'h0000d500, 32'h0000d1fe, 32'h0000d600, 32'h0000d1fe, 32'h0000d700, 
32'h0000d1fe, 32'h0000d800, 32'h0000d1fe, 32'h0000d900, 32'h0000d1fe, 32'h0000da00, 32'h0000d1fe, 32'h0000db00, 32'h0000d1fe, 32'h0000dc00, 32'h0000d1fe, 32'h0000dd00, 32'h0000d1fe, 32'h0000de00, 32'h0000d1fe, 32'h0000df00, 
32'h0000df8d, 32'h0000e000, 32'h0000df8d, 32'h0000e100, 32'h0000df8d, 32'h0000e200, 32'h0000df8d, 32'h0000e300, 32'h0000df8d, 32'h0000e400, 32'h0000df8d, 32'h0000e500, 32'h0000df8d, 32'h0000e600, 32'h0000df8d, 32'h0000e700, 
32'h0000df8d, 32'h0000e800, 32'h0000df8d, 32'h0000e900, 32'h0000df8d, 32'h0000ea00, 32'h0000df8d, 32'h0000eb00, 32'h0000ea8d, 32'h0000ec00, 32'h0000ea8d, 32'h0000ed00, 32'h0000ea8d, 32'h0000ee00, 32'h0000ea8d, 32'h0000ef00, 
32'h0000ea8d, 32'h0000f000, 32'h0000ea8d, 32'h0000f100, 32'h0000ea8d, 32'h0000f200, 32'h0000ea8d, 32'h0000f300, 32'h0000ea8d, 32'h0000f400, 32'h0000ea8d, 32'h0000f500, 32'h0000ea8d, 32'h0000f600, 32'h0000f5c6, 32'h0000f700, 
32'h0000f5c6, 32'h0000f800, 32'h0000f5c6, 32'h0000f900, 32'h0000f5c6, 32'h0000fa00, 32'h0000f5c6, 32'h0000fb00, 32'h0000fae3, 32'h0000fc00, 32'h0000fae3, 32'h0000fd00, 32'h0000fce3, 32'h0000fe00, 32'h0000fce3, 32'h0000ff00 
};

assign slot_freqs={
32'h00000639, 32'h00000000, 32'h00000639, 32'h00000000, 32'h00000639, 32'h00000000, 32'h00000639, 32'h00000000, 32'h00000639, 32'h00000000, 32'h00000639, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 
32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000639, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 
32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 
32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 
32'h0000031c, 32'h0000255a, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 
32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000255a, 32'h00000000, 32'h0000018f, 32'h0000031c, 32'h00000256, 32'h0000018f, 32'h0000031c, 32'h000000c7, 32'h0000031c, 32'h00000000, 
32'h0000031c, 32'h00000000, 32'h0000018f, 32'h00000000, 32'h00000256, 32'h00000000, 32'h0000018e, 32'h00000000, 32'h00000256, 32'h00000000, 32'h00000256, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 
32'h000003e4, 32'h00000000, 32'h00000255, 32'h00000000, 32'h00000255, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 
32'h000003e4, 32'h00000000, 32'h0000031d, 32'h00000256, 32'h0000031d, 32'h00000000, 32'h0000031d, 32'h0000018e, 32'h0000031d, 32'h00000256, 32'h00000256, 32'h000003e4, 32'h00000256, 32'h00000255, 32'h00000256, 32'h00000000, 
32'h00000256, 32'h000000c7, 32'h00000256, 32'h0000031d, 32'h00000256, 32'h00000000, 32'h00000ae5, 32'h000000c7, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h000000c7, 32'h00000ae5, 32'h000003e4, 32'h00000ae5, 32'h0000031d, 
32'h00000ae5, 32'h000000c7, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000256, 32'h00000ae5, 32'h000000c7, 32'h00000ae5, 32'h00000256, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h000000c7, 
32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000572, 32'h00000000, 32'h00000572, 32'h00000000, 32'h00000572, 32'h00000000, 32'h00000572, 32'h00000000, 32'h00000572, 32'h00000000, 
32'h0000088f, 32'h00000000, 32'h0000088f, 32'h00000ae5, 32'h0000088f, 32'h00000000, 32'h0000088f, 32'h00000572, 32'h0000181f, 32'h0000088f, 32'h00000256, 32'h0000181f, 32'h0000031d, 32'h00000256, 32'h00000ae5, 32'h0000031d, 
32'h00000f90, 32'h00000ae5, 32'h000003e4, 32'h00000f90, 32'h0000088f, 32'h00000000, 32'h000003e4, 32'h000003e4, 32'h000004ab, 32'h000003e4, 32'h0000111e, 32'h000004ab, 32'h000007c8, 32'h0000111e, 32'h000003e4, 32'h000007c8, 
32'h00000e02, 32'h000003e4, 32'h0000088f, 32'h00000000, 32'h00000c73, 32'h00000e02, 32'h00000c73, 32'h00000c73, 32'h0000063a, 32'h00000c73, 32'h0000031d, 32'h0000063a, 32'h0000088f, 32'h000000c7, 32'h0000031d, 32'h0000031d, 
32'h0000088f, 32'h000000c7, 32'h0000031d, 32'h0000031d, 32'h0000088f, 32'h00000000, 32'h0000088f, 32'h00000000, 32'h0000088f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 
32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 
32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 
32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h0000181f, 32'h00000000, 32'h00000256, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h00000ae5, 32'h00000000, 
32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 32'h00000ae5, 32'h00000000, 
32'h00000ae5, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 
32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 32'h00000f90, 32'h00000000, 
32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000004ab, 32'h00000000, 32'h000004ab, 32'h00000000, 
32'h000004ab, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 
32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 32'h0000111e, 32'h00000000, 
32'h0000111e, 32'h00000000, 32'h000007c8, 32'h00000000, 32'h000007c8, 32'h00000000, 32'h000007c8, 32'h00000000, 32'h000007c8, 32'h00000000, 32'h000007c8, 32'h00000000, 32'h000007c8, 32'h00000000, 32'h000007c8, 32'h00000000, 
32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h000003e4, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 
32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 32'h00000e02, 32'h00000000, 
32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 
32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 
32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h00000c73, 32'h00000000, 32'h0000063a, 32'h00000000, 
32'h0000063a, 32'h00000000, 32'h0000063a, 32'h00000000, 32'h0000063a, 32'h00000000, 32'h0000063a, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h0000031d, 32'h00000000, 32'h0000031d, 32'h00000000 
};

assign sym_id={
32'h0000000a, 32'h00000000, 32'h0000000a, 32'h00000001, 32'h0000000a, 32'h00000002, 32'h0000000a, 32'h00000003, 32'h0000000a, 32'h00000004, 32'h0000000a, 32'h00000005, 32'h00000020, 32'h00000006, 32'h00000020, 32'h00000007, 
32'h00000020, 32'h00000008, 32'h00000020, 32'h00000009, 32'h00000020, 32'h0000000a, 32'h00000020, 32'h0000000b, 32'h00000020, 32'h0000000c, 32'h00000020, 32'h0000000d, 32'h00000020, 32'h0000000e, 32'h00000020, 32'h0000000f, 
32'h00000020, 32'h00000010, 32'h00000020, 32'h00000011, 32'h00000020, 32'h00000012, 32'h00000020, 32'h00000013, 32'h00000020, 32'h00000014, 32'h00000020, 32'h00000015, 32'h00000020, 32'h00000016, 32'h00000020, 32'h00000017, 
32'h00000020, 32'h00000018, 32'h00000020, 32'h00000019, 32'h00000020, 32'h0000001a, 32'h00000020, 32'h0000001b, 32'h00000020, 32'h0000001c, 32'h00000020, 32'h0000001d, 32'h00000020, 32'h0000001e, 32'h00000020, 32'h0000001f, 
32'h0000002c, 32'h00000020, 32'h00000020, 32'h00000021, 32'h00000020, 32'h00000022, 32'h00000020, 32'h00000023, 32'h00000020, 32'h00000024, 32'h00000020, 32'h00000025, 32'h00000020, 32'h00000026, 32'h00000020, 32'h00000027, 
32'h00000020, 32'h00000028, 32'h00000020, 32'h00000029, 32'h00000020, 32'h0000002a, 32'h00000020, 32'h0000002b, 32'h0000002d, 32'h0000002c, 32'h00000041, 32'h0000002d, 32'h0000002c, 32'h0000002e, 32'h0000002c, 32'h0000002f, 
32'h0000002c, 32'h00000030, 32'h0000002d, 32'h00000031, 32'h00000041, 32'h00000032, 32'h00000043, 32'h00000033, 32'h00000044, 32'h00000034, 32'h00000044, 32'h00000035, 32'h00000045, 32'h00000036, 32'h00000045, 32'h00000037, 
32'h00000045, 32'h00000038, 32'h00000046, 32'h00000039, 32'h00000046, 32'h0000003a, 32'h00000049, 32'h0000003b, 32'h00000049, 32'h0000003c, 32'h00000049, 32'h0000003d, 32'h0000004e, 32'h0000003e, 32'h0000004e, 32'h0000003f, 
32'h0000004e, 32'h00000040, 32'h0000004f, 32'h00000041, 32'h0000004f, 32'h00000042, 32'h0000004f, 32'h00000043, 32'h0000004f, 32'h00000044, 32'h00000052, 32'h00000045, 32'h00000052, 32'h00000046, 32'h00000052, 32'h00000047, 
32'h00000054, 32'h00000048, 32'h00000054, 32'h00000049, 32'h00000054, 32'h0000004a, 32'h00000061, 32'h0000004b, 32'h00000061, 32'h0000004c, 32'h00000061, 32'h0000004d, 32'h00000061, 32'h0000004e, 32'h00000061, 32'h0000004f, 
32'h00000061, 32'h00000050, 32'h00000061, 32'h00000051, 32'h00000061, 32'h00000052, 32'h00000061, 32'h00000053, 32'h00000061, 32'h00000054, 32'h00000061, 32'h00000055, 32'h00000061, 32'h00000056, 32'h00000061, 32'h00000057, 
32'h00000061, 32'h00000058, 32'h00000061, 32'h00000059, 32'h00000061, 32'h0000005a, 32'h00000063, 32'h0000005b, 32'h00000063, 32'h0000005c, 32'h00000063, 32'h0000005d, 32'h00000063, 32'h0000005e, 32'h00000063, 32'h0000005f, 
32'h00000064, 32'h00000060, 32'h00000064, 32'h00000061, 32'h00000064, 32'h00000062, 32'h00000064, 32'h00000063, 32'h00000065, 32'h00000064, 32'h00000066, 32'h00000065, 32'h00000067, 32'h00000066, 32'h00000068, 32'h00000067, 
32'h00000069, 32'h00000068, 32'h0000006b, 32'h00000069, 32'h00000064, 32'h0000006a, 32'h0000006c, 32'h0000006b, 32'h0000006d, 32'h0000006c, 32'h0000006e, 32'h0000006d, 32'h0000006f, 32'h0000006e, 32'h00000070, 32'h0000006f, 
32'h00000072, 32'h00000070, 32'h00000064, 32'h00000071, 32'h00000073, 32'h00000072, 32'h00000074, 32'h00000073, 32'h00000075, 32'h00000074, 32'h00000077, 32'h00000075, 32'h00000064, 32'h00000076, 32'h00000079, 32'h00000077, 
32'h00000064, 32'h00000078, 32'h00000079, 32'h00000079, 32'h00000064, 32'h0000007a, 32'h00000064, 32'h0000007b, 32'h00000064, 32'h0000007c, 32'h00000065, 32'h0000007d, 32'h00000065, 32'h0000007e, 32'h00000065, 32'h0000007f, 
32'h00000065, 32'h00000080, 32'h00000065, 32'h00000081, 32'h00000065, 32'h00000082, 32'h00000065, 32'h00000083, 32'h00000065, 32'h00000084, 32'h00000065, 32'h00000085, 32'h00000065, 32'h00000086, 32'h00000065, 32'h00000087, 
32'h00000065, 32'h00000088, 32'h00000065, 32'h00000089, 32'h00000065, 32'h0000008a, 32'h00000065, 32'h0000008b, 32'h00000065, 32'h0000008c, 32'h00000065, 32'h0000008d, 32'h00000065, 32'h0000008e, 32'h00000065, 32'h0000008f, 
32'h00000065, 32'h00000090, 32'h00000065, 32'h00000091, 32'h00000065, 32'h00000092, 32'h00000065, 32'h00000093, 32'h00000066, 32'h00000094, 32'h00000067, 32'h00000095, 32'h00000067, 32'h00000096, 32'h00000068, 32'h00000097, 
32'h00000068, 32'h00000098, 32'h00000068, 32'h00000099, 32'h00000068, 32'h0000009a, 32'h00000068, 32'h0000009b, 32'h00000068, 32'h0000009c, 32'h00000068, 32'h0000009d, 32'h00000068, 32'h0000009e, 32'h00000068, 32'h0000009f, 
32'h00000068, 32'h000000a0, 32'h00000069, 32'h000000a1, 32'h00000069, 32'h000000a2, 32'h00000069, 32'h000000a3, 32'h00000069, 32'h000000a4, 32'h00000069, 32'h000000a5, 32'h00000069, 32'h000000a6, 32'h00000069, 32'h000000a7, 
32'h00000069, 32'h000000a8, 32'h00000069, 32'h000000a9, 32'h00000069, 32'h000000aa, 32'h00000069, 32'h000000ab, 32'h00000069, 32'h000000ac, 32'h00000069, 32'h000000ad, 32'h00000069, 32'h000000ae, 32'h00000069, 32'h000000af, 
32'h0000006b, 32'h000000b0, 32'h0000006b, 32'h000000b1, 32'h0000006b, 32'h000000b2, 32'h0000006c, 32'h000000b3, 32'h0000006c, 32'h000000b4, 32'h0000006c, 32'h000000b5, 32'h0000006d, 32'h000000b6, 32'h0000006d, 32'h000000b7, 
32'h0000006d, 32'h000000b8, 32'h0000006e, 32'h000000b9, 32'h0000006e, 32'h000000ba, 32'h0000006e, 32'h000000bb, 32'h0000006e, 32'h000000bc, 32'h0000006e, 32'h000000bd, 32'h0000006e, 32'h000000be, 32'h0000006e, 32'h000000bf, 
32'h0000006e, 32'h000000c0, 32'h0000006e, 32'h000000c1, 32'h0000006e, 32'h000000c2, 32'h0000006e, 32'h000000c3, 32'h0000006e, 32'h000000c4, 32'h0000006e, 32'h000000c5, 32'h0000006e, 32'h000000c6, 32'h0000006e, 32'h000000c7, 
32'h0000006e, 32'h000000c8, 32'h0000006f, 32'h000000c9, 32'h0000006f, 32'h000000ca, 32'h0000006f, 32'h000000cb, 32'h0000006f, 32'h000000cc, 32'h0000006f, 32'h000000cd, 32'h0000006f, 32'h000000ce, 32'h0000006f, 32'h000000cf, 
32'h00000070, 32'h000000d0, 32'h00000070, 32'h000000d1, 32'h00000070, 32'h000000d2, 32'h00000072, 32'h000000d3, 32'h00000072, 32'h000000d4, 32'h00000072, 32'h000000d5, 32'h00000072, 32'h000000d6, 32'h00000072, 32'h000000d7, 
32'h00000072, 32'h000000d8, 32'h00000072, 32'h000000d9, 32'h00000072, 32'h000000da, 32'h00000072, 32'h000000db, 32'h00000072, 32'h000000dc, 32'h00000072, 32'h000000dd, 32'h00000072, 32'h000000de, 32'h00000072, 32'h000000df, 
32'h00000073, 32'h000000e0, 32'h00000073, 32'h000000e1, 32'h00000073, 32'h000000e2, 32'h00000073, 32'h000000e3, 32'h00000073, 32'h000000e4, 32'h00000073, 32'h000000e5, 32'h00000073, 32'h000000e6, 32'h00000073, 32'h000000e7, 
32'h00000073, 32'h000000e8, 32'h00000073, 32'h000000e9, 32'h00000073, 32'h000000ea, 32'h00000073, 32'h000000eb, 32'h00000074, 32'h000000ec, 32'h00000074, 32'h000000ed, 32'h00000074, 32'h000000ee, 32'h00000074, 32'h000000ef, 
32'h00000074, 32'h000000f0, 32'h00000074, 32'h000000f1, 32'h00000074, 32'h000000f2, 32'h00000074, 32'h000000f3, 32'h00000074, 32'h000000f4, 32'h00000074, 32'h000000f5, 32'h00000074, 32'h000000f6, 32'h00000075, 32'h000000f7, 
32'h00000075, 32'h000000f8, 32'h00000075, 32'h000000f9, 32'h00000075, 32'h000000fa, 32'h00000075, 32'h000000fb, 32'h00000077, 32'h000000fc, 32'h00000077, 32'h000000fd, 32'h00000079, 32'h000000fe, 32'h00000079, 32'h000000ff 
};
// End of Computer Generated tables:


endmodule


